
module aes_improve_critical_paths
(
  done,
  text_out,
  text_in_r,
  sa00,
  sa01,
  sa02,
  sa03,
  sa10,
  sa11,
  sa12,
  sa13,
  sa20,
  sa21,
  sa22,
  sa23,
  sa30,
  sa31,
  sa32,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33,
  sa33
);

  assign Cond42 = sa00;
  assign ld_r = Cond42;
  assign Cond34 = sa01;
  assign ld_r = Cond34;
  assign Cond26 = sa02;
  assign ld_r = Cond26;
  assign Cond18 = sa03;
  assign ld_r = Cond18;
  assign Cond40 = sa10;
  assign ld_r = Cond40;
  assign Cond32 = sa11;
  assign ld_r = Cond32;
  assign Cond24 = sa12;
  assign ld_r = Cond24;
  assign Cond16 = sa13;
  assign ld_r = Cond16;
  assign Cond38 = sa20;
  assign ld_r = Cond38;
  assign Cond30 = sa21;
  assign ld_r = Cond30;
  assign Cond22 = sa22;
  assign ld_r = Cond22;
  assign Cond14 = sa23;
  assign ld_r = Cond14;
  assign Cond36 = sa30;
  assign ld_r = Cond36;
  assign Cond28 = sa31;
  assign ld_r = Cond28;
  assign Cond20 = sa32;
  assign ld_r = Cond20;
  assign Cond12 = sa33;
  assign ld_r = Cond12;

endmodule
